LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all;

ENTITY afficheur7segment IS
    PORT (ck, rst: IN STD_LOGIC;
           q : out STD_LOGIC);
END afficheur7segment;

ARCHITECTURE program OF afficheur7segment IS
BEGIN 
        
     
END program;